
`timescale 1ns / 1ps
module dromi_16x512 #(
    parameter    ADDR_WIDTH     =   9,
    parameter    DATA_WIDTH     =   16
) (
    input   wire                        clk,
    input   wire                        rst,
    input   wire                        clk_en,

    input   wire    [ADDR_WIDTH-1:0]    addr,
    output  reg     [DATA_WIDTH-1:0]    rd_data
);

always@(posedge clk or posedge rst) begin
    if (rst) begin
		rd_data <= 0;
	end
	else begin
		if(clk_en) begin
			case (addr)
				0	: begin rd_data <= 16'h0000; end
				1	: begin rd_data <= 16'hff9b; end
				2	: begin rd_data <= 16'hff37; end
				3	: begin rd_data <= 16'hfed2; end
				4	: begin rd_data <= 16'hfe6e; end
				5	: begin rd_data <= 16'hfe09; end
				6	: begin rd_data <= 16'hfda5; end
				7	: begin rd_data <= 16'hfd40; end
				8	: begin rd_data <= 16'hfcdc; end
				9	: begin rd_data <= 16'hfc78; end
				10	: begin rd_data <= 16'hfc13; end
				11	: begin rd_data <= 16'hfbaf; end
				12	: begin rd_data <= 16'hfb4b; end
				13	: begin rd_data <= 16'hfae6; end
				14	: begin rd_data <= 16'hfa82; end
				15	: begin rd_data <= 16'hfa1e; end
				16	: begin rd_data <= 16'hf9ba; end
				17	: begin rd_data <= 16'hf956; end
				18	: begin rd_data <= 16'hf8f2; end
				19	: begin rd_data <= 16'hf88e; end
				20	: begin rd_data <= 16'hf82a; end
				21	: begin rd_data <= 16'hf7c7; end
				22	: begin rd_data <= 16'hf763; end
				23	: begin rd_data <= 16'hf6ff; end
				24	: begin rd_data <= 16'hf69c; end
				25	: begin rd_data <= 16'hf639; end
				26	: begin rd_data <= 16'hf5d5; end
				27	: begin rd_data <= 16'hf572; end
				28	: begin rd_data <= 16'hf50f; end
				29	: begin rd_data <= 16'hf4ac; end
				30	: begin rd_data <= 16'hf449; end
				31	: begin rd_data <= 16'hf3e6; end
				32	: begin rd_data <= 16'hf384; end
				33	: begin rd_data <= 16'hf321; end
				34	: begin rd_data <= 16'hf2bf; end
				35	: begin rd_data <= 16'hf25c; end
				36	: begin rd_data <= 16'hf1fa; end
				37	: begin rd_data <= 16'hf198; end
				38	: begin rd_data <= 16'hf136; end
				39	: begin rd_data <= 16'hf0d5; end
				40	: begin rd_data <= 16'hf073; end
				41	: begin rd_data <= 16'hf012; end
				42	: begin rd_data <= 16'hefb0; end
				43	: begin rd_data <= 16'hef4f; end
				44	: begin rd_data <= 16'heeee; end
				45	: begin rd_data <= 16'hee8d; end
				46	: begin rd_data <= 16'hee2d; end
				47	: begin rd_data <= 16'hedcc; end
				48	: begin rd_data <= 16'hed6c; end
				49	: begin rd_data <= 16'hed0c; end
				50	: begin rd_data <= 16'hecac; end
				51	: begin rd_data <= 16'hec4c; end
				52	: begin rd_data <= 16'hebed; end
				53	: begin rd_data <= 16'heb8d; end
				54	: begin rd_data <= 16'heb2e; end
				55	: begin rd_data <= 16'heacf; end
				56	: begin rd_data <= 16'hea70; end
				57	: begin rd_data <= 16'hea12; end
				58	: begin rd_data <= 16'he9b4; end
				59	: begin rd_data <= 16'he955; end
				60	: begin rd_data <= 16'he8f7; end
				61	: begin rd_data <= 16'he89a; end
				62	: begin rd_data <= 16'he83c; end
				63	: begin rd_data <= 16'he7df; end
				64	: begin rd_data <= 16'he782; end
				65	: begin rd_data <= 16'he725; end
				66	: begin rd_data <= 16'he6c9; end
				67	: begin rd_data <= 16'he66d; end
				68	: begin rd_data <= 16'he611; end
				69	: begin rd_data <= 16'he5b5; end
				70	: begin rd_data <= 16'he559; end
				71	: begin rd_data <= 16'he4fe; end
				72	: begin rd_data <= 16'he4a3; end
				73	: begin rd_data <= 16'he448; end
				74	: begin rd_data <= 16'he3ee; end
				75	: begin rd_data <= 16'he394; end
				76	: begin rd_data <= 16'he33a; end
				77	: begin rd_data <= 16'he2e0; end
				78	: begin rd_data <= 16'he287; end
				79	: begin rd_data <= 16'he22d; end
				80	: begin rd_data <= 16'he1d5; end
				81	: begin rd_data <= 16'he17c; end
				82	: begin rd_data <= 16'he124; end
				83	: begin rd_data <= 16'he0cc; end
				84	: begin rd_data <= 16'he074; end
				85	: begin rd_data <= 16'he01d; end
				86	: begin rd_data <= 16'hdfc6; end
				87	: begin rd_data <= 16'hdf6f; end
				88	: begin rd_data <= 16'hdf19; end
				89	: begin rd_data <= 16'hdec3; end
				90	: begin rd_data <= 16'hde6d; end
				91	: begin rd_data <= 16'hde18; end
				92	: begin rd_data <= 16'hddc3; end
				93	: begin rd_data <= 16'hdd6e; end
				94	: begin rd_data <= 16'hdd19; end
				95	: begin rd_data <= 16'hdcc5; end
				96	: begin rd_data <= 16'hdc72; end
				97	: begin rd_data <= 16'hdc1e; end
				98	: begin rd_data <= 16'hdbcb; end
				99	: begin rd_data <= 16'hdb78; end
				100	: begin rd_data <= 16'hdb26; end
				101	: begin rd_data <= 16'hdad4; end
				102	: begin rd_data <= 16'hda82; end
				103	: begin rd_data <= 16'hda31; end
				104	: begin rd_data <= 16'hd9e0; end
				105	: begin rd_data <= 16'hd98f; end
				106	: begin rd_data <= 16'hd93f; end
				107	: begin rd_data <= 16'hd8ef; end
				108	: begin rd_data <= 16'hd8a0; end
				109	: begin rd_data <= 16'hd851; end
				110	: begin rd_data <= 16'hd802; end
				111	: begin rd_data <= 16'hd7b4; end
				112	: begin rd_data <= 16'hd766; end
				113	: begin rd_data <= 16'hd719; end
				114	: begin rd_data <= 16'hd6cb; end
				115	: begin rd_data <= 16'hd67f; end
				116	: begin rd_data <= 16'hd632; end
				117	: begin rd_data <= 16'hd5e6; end
				118	: begin rd_data <= 16'hd59b; end
				119	: begin rd_data <= 16'hd550; end
				120	: begin rd_data <= 16'hd505; end
				121	: begin rd_data <= 16'hd4bb; end
				122	: begin rd_data <= 16'hd471; end
				123	: begin rd_data <= 16'hd428; end
				124	: begin rd_data <= 16'hd3df; end
				125	: begin rd_data <= 16'hd396; end
				126	: begin rd_data <= 16'hd34e; end
				127	: begin rd_data <= 16'hd306; end
				128	: begin rd_data <= 16'hd2bf; end
				129	: begin rd_data <= 16'hd278; end
				130	: begin rd_data <= 16'hd231; end
				131	: begin rd_data <= 16'hd1eb; end
				132	: begin rd_data <= 16'hd1a6; end
				133	: begin rd_data <= 16'hd161; end
				134	: begin rd_data <= 16'hd11c; end
				135	: begin rd_data <= 16'hd0d8; end
				136	: begin rd_data <= 16'hd094; end
				137	: begin rd_data <= 16'hd051; end
				138	: begin rd_data <= 16'hd00e; end
				139	: begin rd_data <= 16'hcfcc; end
				140	: begin rd_data <= 16'hcf8a; end
				141	: begin rd_data <= 16'hcf48; end
				142	: begin rd_data <= 16'hcf07; end
				143	: begin rd_data <= 16'hcec7; end
				144	: begin rd_data <= 16'hce87; end
				145	: begin rd_data <= 16'hce47; end
				146	: begin rd_data <= 16'hce08; end
				147	: begin rd_data <= 16'hcdca; end
				148	: begin rd_data <= 16'hcd8c; end
				149	: begin rd_data <= 16'hcd4e; end
				150	: begin rd_data <= 16'hcd11; end
				151	: begin rd_data <= 16'hccd4; end
				152	: begin rd_data <= 16'hcc98; end
				153	: begin rd_data <= 16'hcc5d; end
				154	: begin rd_data <= 16'hcc21; end
				155	: begin rd_data <= 16'hcbe7; end
				156	: begin rd_data <= 16'hcbad; end
				157	: begin rd_data <= 16'hcb73; end
				158	: begin rd_data <= 16'hcb3a; end
				159	: begin rd_data <= 16'hcb01; end
				160	: begin rd_data <= 16'hcac9; end
				161	: begin rd_data <= 16'hca92; end
				162	: begin rd_data <= 16'hca5b; end
				163	: begin rd_data <= 16'hca24; end
				164	: begin rd_data <= 16'hc9ee; end
				165	: begin rd_data <= 16'hc9b8; end
				166	: begin rd_data <= 16'hc983; end
				167	: begin rd_data <= 16'hc94f; end
				168	: begin rd_data <= 16'hc91b; end
				169	: begin rd_data <= 16'hc8e8; end
				170	: begin rd_data <= 16'hc8b5; end
				171	: begin rd_data <= 16'hc882; end
				172	: begin rd_data <= 16'hc850; end
				173	: begin rd_data <= 16'hc81f; end
				174	: begin rd_data <= 16'hc7ee; end
				175	: begin rd_data <= 16'hc7be; end
				176	: begin rd_data <= 16'hc78f; end
				177	: begin rd_data <= 16'hc75f; end
				178	: begin rd_data <= 16'hc731; end
				179	: begin rd_data <= 16'hc703; end
				180	: begin rd_data <= 16'hc6d5; end
				181	: begin rd_data <= 16'hc6a8; end
				182	: begin rd_data <= 16'hc67c; end
				183	: begin rd_data <= 16'hc650; end
				184	: begin rd_data <= 16'hc625; end
				185	: begin rd_data <= 16'hc5fa; end
				186	: begin rd_data <= 16'hc5d0; end
				187	: begin rd_data <= 16'hc5a7; end
				188	: begin rd_data <= 16'hc57e; end
				189	: begin rd_data <= 16'hc555; end
				190	: begin rd_data <= 16'hc52d; end
				191	: begin rd_data <= 16'hc506; end
				192	: begin rd_data <= 16'hc4df; end
				193	: begin rd_data <= 16'hc4b9; end
				194	: begin rd_data <= 16'hc493; end
				195	: begin rd_data <= 16'hc46e; end
				196	: begin rd_data <= 16'hc44a; end
				197	: begin rd_data <= 16'hc426; end
				198	: begin rd_data <= 16'hc403; end
				199	: begin rd_data <= 16'hc3e0; end
				200	: begin rd_data <= 16'hc3be; end
				201	: begin rd_data <= 16'hc39c; end
				202	: begin rd_data <= 16'hc37b; end
				203	: begin rd_data <= 16'hc35b; end
				204	: begin rd_data <= 16'hc33b; end
				205	: begin rd_data <= 16'hc31c; end
				206	: begin rd_data <= 16'hc2fd; end
				207	: begin rd_data <= 16'hc2df; end
				208	: begin rd_data <= 16'hc2c1; end
				209	: begin rd_data <= 16'hc2a5; end
				210	: begin rd_data <= 16'hc288; end
				211	: begin rd_data <= 16'hc26d; end
				212	: begin rd_data <= 16'hc251; end
				213	: begin rd_data <= 16'hc237; end
				214	: begin rd_data <= 16'hc21d; end
				215	: begin rd_data <= 16'hc204; end
				216	: begin rd_data <= 16'hc1eb; end
				217	: begin rd_data <= 16'hc1d3; end
				218	: begin rd_data <= 16'hc1bb; end
				219	: begin rd_data <= 16'hc1a4; end
				220	: begin rd_data <= 16'hc18e; end
				221	: begin rd_data <= 16'hc178; end
				222	: begin rd_data <= 16'hc163; end
				223	: begin rd_data <= 16'hc14f; end
				224	: begin rd_data <= 16'hc13b; end
				225	: begin rd_data <= 16'hc128; end
				226	: begin rd_data <= 16'hc115; end
				227	: begin rd_data <= 16'hc103; end
				228	: begin rd_data <= 16'hc0f1; end
				229	: begin rd_data <= 16'hc0e0; end
				230	: begin rd_data <= 16'hc0d0; end
				231	: begin rd_data <= 16'hc0c0; end
				232	: begin rd_data <= 16'hc0b1; end
				233	: begin rd_data <= 16'hc0a3; end
				234	: begin rd_data <= 16'hc095; end
				235	: begin rd_data <= 16'hc088; end
				236	: begin rd_data <= 16'hc07b; end
				237	: begin rd_data <= 16'hc06f; end
				238	: begin rd_data <= 16'hc064; end
				239	: begin rd_data <= 16'hc059; end
				240	: begin rd_data <= 16'hc04f; end
				241	: begin rd_data <= 16'hc045; end
				242	: begin rd_data <= 16'hc03c; end
				243	: begin rd_data <= 16'hc034; end
				244	: begin rd_data <= 16'hc02c; end
				245	: begin rd_data <= 16'hc025; end
				246	: begin rd_data <= 16'hc01f; end
				247	: begin rd_data <= 16'hc019; end
				248	: begin rd_data <= 16'hc014; end
				249	: begin rd_data <= 16'hc00f; end
				250	: begin rd_data <= 16'hc00b; end
				251	: begin rd_data <= 16'hc008; end
				252	: begin rd_data <= 16'hc005; end
				253	: begin rd_data <= 16'hc003; end
				254	: begin rd_data <= 16'hc001; end
				255	: begin rd_data <= 16'hc000; end
				256	: begin rd_data <= 16'hc000; end
				257	: begin rd_data <= 16'hc000; end
				258	: begin rd_data <= 16'hc001; end
				259	: begin rd_data <= 16'hc003; end
				260	: begin rd_data <= 16'hc005; end
				261	: begin rd_data <= 16'hc008; end
				262	: begin rd_data <= 16'hc00b; end
				263	: begin rd_data <= 16'hc00f; end
				264	: begin rd_data <= 16'hc014; end
				265	: begin rd_data <= 16'hc019; end
				266	: begin rd_data <= 16'hc01f; end
				267	: begin rd_data <= 16'hc025; end
				268	: begin rd_data <= 16'hc02c; end
				269	: begin rd_data <= 16'hc034; end
				270	: begin rd_data <= 16'hc03c; end
				271	: begin rd_data <= 16'hc045; end
				272	: begin rd_data <= 16'hc04f; end
				273	: begin rd_data <= 16'hc059; end
				274	: begin rd_data <= 16'hc064; end
				275	: begin rd_data <= 16'hc06f; end
				276	: begin rd_data <= 16'hc07b; end
				277	: begin rd_data <= 16'hc088; end
				278	: begin rd_data <= 16'hc095; end
				279	: begin rd_data <= 16'hc0a3; end
				280	: begin rd_data <= 16'hc0b1; end
				281	: begin rd_data <= 16'hc0c0; end
				282	: begin rd_data <= 16'hc0d0; end
				283	: begin rd_data <= 16'hc0e0; end
				284	: begin rd_data <= 16'hc0f1; end
				285	: begin rd_data <= 16'hc103; end
				286	: begin rd_data <= 16'hc115; end
				287	: begin rd_data <= 16'hc128; end
				288	: begin rd_data <= 16'hc13b; end
				289	: begin rd_data <= 16'hc14f; end
				290	: begin rd_data <= 16'hc163; end
				291	: begin rd_data <= 16'hc178; end
				292	: begin rd_data <= 16'hc18e; end
				293	: begin rd_data <= 16'hc1a4; end
				294	: begin rd_data <= 16'hc1bb; end
				295	: begin rd_data <= 16'hc1d3; end
				296	: begin rd_data <= 16'hc1eb; end
				297	: begin rd_data <= 16'hc204; end
				298	: begin rd_data <= 16'hc21d; end
				299	: begin rd_data <= 16'hc237; end
				300	: begin rd_data <= 16'hc251; end
				301	: begin rd_data <= 16'hc26d; end
				302	: begin rd_data <= 16'hc288; end
				303	: begin rd_data <= 16'hc2a5; end
				304	: begin rd_data <= 16'hc2c1; end
				305	: begin rd_data <= 16'hc2df; end
				306	: begin rd_data <= 16'hc2fd; end
				307	: begin rd_data <= 16'hc31c; end
				308	: begin rd_data <= 16'hc33b; end
				309	: begin rd_data <= 16'hc35b; end
				310	: begin rd_data <= 16'hc37b; end
				311	: begin rd_data <= 16'hc39c; end
				312	: begin rd_data <= 16'hc3be; end
				313	: begin rd_data <= 16'hc3e0; end
				314	: begin rd_data <= 16'hc403; end
				315	: begin rd_data <= 16'hc426; end
				316	: begin rd_data <= 16'hc44a; end
				317	: begin rd_data <= 16'hc46e; end
				318	: begin rd_data <= 16'hc493; end
				319	: begin rd_data <= 16'hc4b9; end
				320	: begin rd_data <= 16'hc4df; end
				321	: begin rd_data <= 16'hc506; end
				322	: begin rd_data <= 16'hc52d; end
				323	: begin rd_data <= 16'hc555; end
				324	: begin rd_data <= 16'hc57e; end
				325	: begin rd_data <= 16'hc5a7; end
				326	: begin rd_data <= 16'hc5d0; end
				327	: begin rd_data <= 16'hc5fa; end
				328	: begin rd_data <= 16'hc625; end
				329	: begin rd_data <= 16'hc650; end
				330	: begin rd_data <= 16'hc67c; end
				331	: begin rd_data <= 16'hc6a8; end
				332	: begin rd_data <= 16'hc6d5; end
				333	: begin rd_data <= 16'hc703; end
				334	: begin rd_data <= 16'hc731; end
				335	: begin rd_data <= 16'hc75f; end
				336	: begin rd_data <= 16'hc78f; end
				337	: begin rd_data <= 16'hc7be; end
				338	: begin rd_data <= 16'hc7ee; end
				339	: begin rd_data <= 16'hc81f; end
				340	: begin rd_data <= 16'hc850; end
				341	: begin rd_data <= 16'hc882; end
				342	: begin rd_data <= 16'hc8b5; end
				343	: begin rd_data <= 16'hc8e8; end
				344	: begin rd_data <= 16'hc91b; end
				345	: begin rd_data <= 16'hc94f; end
				346	: begin rd_data <= 16'hc983; end
				347	: begin rd_data <= 16'hc9b8; end
				348	: begin rd_data <= 16'hc9ee; end
				349	: begin rd_data <= 16'hca24; end
				350	: begin rd_data <= 16'hca5b; end
				351	: begin rd_data <= 16'hca92; end
				352	: begin rd_data <= 16'hcac9; end
				353	: begin rd_data <= 16'hcb01; end
				354	: begin rd_data <= 16'hcb3a; end
				355	: begin rd_data <= 16'hcb73; end
				356	: begin rd_data <= 16'hcbad; end
				357	: begin rd_data <= 16'hcbe7; end
				358	: begin rd_data <= 16'hcc21; end
				359	: begin rd_data <= 16'hcc5d; end
				360	: begin rd_data <= 16'hcc98; end
				361	: begin rd_data <= 16'hccd4; end
				362	: begin rd_data <= 16'hcd11; end
				363	: begin rd_data <= 16'hcd4e; end
				364	: begin rd_data <= 16'hcd8c; end
				365	: begin rd_data <= 16'hcdca; end
				366	: begin rd_data <= 16'hce08; end
				367	: begin rd_data <= 16'hce47; end
				368	: begin rd_data <= 16'hce87; end
				369	: begin rd_data <= 16'hcec7; end
				370	: begin rd_data <= 16'hcf07; end
				371	: begin rd_data <= 16'hcf48; end
				372	: begin rd_data <= 16'hcf8a; end
				373	: begin rd_data <= 16'hcfcc; end
				374	: begin rd_data <= 16'hd00e; end
				375	: begin rd_data <= 16'hd051; end
				376	: begin rd_data <= 16'hd094; end
				377	: begin rd_data <= 16'hd0d8; end
				378	: begin rd_data <= 16'hd11c; end
				379	: begin rd_data <= 16'hd161; end
				380	: begin rd_data <= 16'hd1a6; end
				381	: begin rd_data <= 16'hd1eb; end
				382	: begin rd_data <= 16'hd231; end
				383	: begin rd_data <= 16'hd278; end
				384	: begin rd_data <= 16'hd2bf; end
				385	: begin rd_data <= 16'hd306; end
				386	: begin rd_data <= 16'hd34e; end
				387	: begin rd_data <= 16'hd396; end
				388	: begin rd_data <= 16'hd3df; end
				389	: begin rd_data <= 16'hd428; end
				390	: begin rd_data <= 16'hd471; end
				391	: begin rd_data <= 16'hd4bb; end
				392	: begin rd_data <= 16'hd505; end
				393	: begin rd_data <= 16'hd550; end
				394	: begin rd_data <= 16'hd59b; end
				395	: begin rd_data <= 16'hd5e6; end
				396	: begin rd_data <= 16'hd632; end
				397	: begin rd_data <= 16'hd67f; end
				398	: begin rd_data <= 16'hd6cb; end
				399	: begin rd_data <= 16'hd719; end
				400	: begin rd_data <= 16'hd766; end
				401	: begin rd_data <= 16'hd7b4; end
				402	: begin rd_data <= 16'hd802; end
				403	: begin rd_data <= 16'hd851; end
				404	: begin rd_data <= 16'hd8a0; end
				405	: begin rd_data <= 16'hd8ef; end
				406	: begin rd_data <= 16'hd93f; end
				407	: begin rd_data <= 16'hd98f; end
				408	: begin rd_data <= 16'hd9e0; end
				409	: begin rd_data <= 16'hda31; end
				410	: begin rd_data <= 16'hda82; end
				411	: begin rd_data <= 16'hdad4; end
				412	: begin rd_data <= 16'hdb26; end
				413	: begin rd_data <= 16'hdb78; end
				414	: begin rd_data <= 16'hdbcb; end
				415	: begin rd_data <= 16'hdc1e; end
				416	: begin rd_data <= 16'hdc72; end
				417	: begin rd_data <= 16'hdcc5; end
				418	: begin rd_data <= 16'hdd19; end
				419	: begin rd_data <= 16'hdd6e; end
				420	: begin rd_data <= 16'hddc3; end
				421	: begin rd_data <= 16'hde18; end
				422	: begin rd_data <= 16'hde6d; end
				423	: begin rd_data <= 16'hdec3; end
				424	: begin rd_data <= 16'hdf19; end
				425	: begin rd_data <= 16'hdf6f; end
				426	: begin rd_data <= 16'hdfc6; end
				427	: begin rd_data <= 16'he01d; end
				428	: begin rd_data <= 16'he074; end
				429	: begin rd_data <= 16'he0cc; end
				430	: begin rd_data <= 16'he124; end
				431	: begin rd_data <= 16'he17c; end
				432	: begin rd_data <= 16'he1d5; end
				433	: begin rd_data <= 16'he22d; end
				434	: begin rd_data <= 16'he287; end
				435	: begin rd_data <= 16'he2e0; end
				436	: begin rd_data <= 16'he33a; end
				437	: begin rd_data <= 16'he394; end
				438	: begin rd_data <= 16'he3ee; end
				439	: begin rd_data <= 16'he448; end
				440	: begin rd_data <= 16'he4a3; end
				441	: begin rd_data <= 16'he4fe; end
				442	: begin rd_data <= 16'he559; end
				443	: begin rd_data <= 16'he5b5; end
				444	: begin rd_data <= 16'he611; end
				445	: begin rd_data <= 16'he66d; end
				446	: begin rd_data <= 16'he6c9; end
				447	: begin rd_data <= 16'he725; end
				448	: begin rd_data <= 16'he782; end
				449	: begin rd_data <= 16'he7df; end
				450	: begin rd_data <= 16'he83c; end
				451	: begin rd_data <= 16'he89a; end
				452	: begin rd_data <= 16'he8f7; end
				453	: begin rd_data <= 16'he955; end
				454	: begin rd_data <= 16'he9b4; end
				455	: begin rd_data <= 16'hea12; end
				456	: begin rd_data <= 16'hea70; end
				457	: begin rd_data <= 16'heacf; end
				458	: begin rd_data <= 16'heb2e; end
				459	: begin rd_data <= 16'heb8d; end
				460	: begin rd_data <= 16'hebed; end
				461	: begin rd_data <= 16'hec4c; end
				462	: begin rd_data <= 16'hecac; end
				463	: begin rd_data <= 16'hed0c; end
				464	: begin rd_data <= 16'hed6c; end
				465	: begin rd_data <= 16'hedcc; end
				466	: begin rd_data <= 16'hee2d; end
				467	: begin rd_data <= 16'hee8d; end
				468	: begin rd_data <= 16'heeee; end
				469	: begin rd_data <= 16'hef4f; end
				470	: begin rd_data <= 16'hefb0; end
				471	: begin rd_data <= 16'hf012; end
				472	: begin rd_data <= 16'hf073; end
				473	: begin rd_data <= 16'hf0d5; end
				474	: begin rd_data <= 16'hf136; end
				475	: begin rd_data <= 16'hf198; end
				476	: begin rd_data <= 16'hf1fa; end
				477	: begin rd_data <= 16'hf25c; end
				478	: begin rd_data <= 16'hf2bf; end
				479	: begin rd_data <= 16'hf321; end
				480	: begin rd_data <= 16'hf384; end
				481	: begin rd_data <= 16'hf3e6; end
				482	: begin rd_data <= 16'hf449; end
				483	: begin rd_data <= 16'hf4ac; end
				484	: begin rd_data <= 16'hf50f; end
				485	: begin rd_data <= 16'hf572; end
				486	: begin rd_data <= 16'hf5d5; end
				487	: begin rd_data <= 16'hf639; end
				488	: begin rd_data <= 16'hf69c; end
				489	: begin rd_data <= 16'hf6ff; end
				490	: begin rd_data <= 16'hf763; end
				491	: begin rd_data <= 16'hf7c7; end
				492	: begin rd_data <= 16'hf82a; end
				493	: begin rd_data <= 16'hf88e; end
				494	: begin rd_data <= 16'hf8f2; end
				495	: begin rd_data <= 16'hf956; end
				496	: begin rd_data <= 16'hf9ba; end
				497	: begin rd_data <= 16'hfa1e; end
				498	: begin rd_data <= 16'hfa82; end
				499	: begin rd_data <= 16'hfae6; end
				500	: begin rd_data <= 16'hfb4b; end
				501	: begin rd_data <= 16'hfbaf; end
				502	: begin rd_data <= 16'hfc13; end
				503	: begin rd_data <= 16'hfc78; end
				504	: begin rd_data <= 16'hfcdc; end
				505	: begin rd_data <= 16'hfd40; end
				506	: begin rd_data <= 16'hfda5; end
				507	: begin rd_data <= 16'hfe09; end
				508	: begin rd_data <= 16'hfe6e; end
				509	: begin rd_data <= 16'hfed2; end
				510	: begin rd_data <= 16'hff37; end
				511	: begin rd_data <= 16'hff9b; end
				default : begin rd_data <= 0; end
			endcase
		end
		else begin
			rd_data <= rd_data;
		end
	end
end

endmodule
