
`timescale 1ns / 1ps
module dromr_16x512 #(
    parameter    ADDR_WIDTH     =   9,
    parameter    DATA_WIDTH     =   16
) (
    input   wire                        clk,
    input   wire                        rst,
    input   wire                        clk_en,

    input   wire    [ADDR_WIDTH-1:0]    addr,
    output  reg     [DATA_WIDTH-1:0]    rd_data
);

always@(posedge clk or posedge rst) begin
    if (rst) begin
		rd_data <= 0;
	end
	else begin
		if(clk_en) begin
			case (addr)
				0	: begin rd_data <= 16'h4000; end
				1	: begin rd_data <= 16'h4000; end
				2	: begin rd_data <= 16'h3fff; end
				3	: begin rd_data <= 16'h3ffd; end
				4	: begin rd_data <= 16'h3ffb; end
				5	: begin rd_data <= 16'h3ff8; end
				6	: begin rd_data <= 16'h3ff5; end
				7	: begin rd_data <= 16'h3ff1; end
				8	: begin rd_data <= 16'h3fec; end
				9	: begin rd_data <= 16'h3fe7; end
				10	: begin rd_data <= 16'h3fe1; end
				11	: begin rd_data <= 16'h3fdb; end
				12	: begin rd_data <= 16'h3fd4; end
				13	: begin rd_data <= 16'h3fcc; end
				14	: begin rd_data <= 16'h3fc4; end
				15	: begin rd_data <= 16'h3fbb; end
				16	: begin rd_data <= 16'h3fb1; end
				17	: begin rd_data <= 16'h3fa7; end
				18	: begin rd_data <= 16'h3f9c; end
				19	: begin rd_data <= 16'h3f91; end
				20	: begin rd_data <= 16'h3f85; end
				21	: begin rd_data <= 16'h3f78; end
				22	: begin rd_data <= 16'h3f6b; end
				23	: begin rd_data <= 16'h3f5d; end
				24	: begin rd_data <= 16'h3f4f; end
				25	: begin rd_data <= 16'h3f40; end
				26	: begin rd_data <= 16'h3f30; end
				27	: begin rd_data <= 16'h3f20; end
				28	: begin rd_data <= 16'h3f0f; end
				29	: begin rd_data <= 16'h3efd; end
				30	: begin rd_data <= 16'h3eeb; end
				31	: begin rd_data <= 16'h3ed8; end
				32	: begin rd_data <= 16'h3ec5; end
				33	: begin rd_data <= 16'h3eb1; end
				34	: begin rd_data <= 16'h3e9d; end
				35	: begin rd_data <= 16'h3e88; end
				36	: begin rd_data <= 16'h3e72; end
				37	: begin rd_data <= 16'h3e5c; end
				38	: begin rd_data <= 16'h3e45; end
				39	: begin rd_data <= 16'h3e2d; end
				40	: begin rd_data <= 16'h3e15; end
				41	: begin rd_data <= 16'h3dfc; end
				42	: begin rd_data <= 16'h3de3; end
				43	: begin rd_data <= 16'h3dc9; end
				44	: begin rd_data <= 16'h3daf; end
				45	: begin rd_data <= 16'h3d93; end
				46	: begin rd_data <= 16'h3d78; end
				47	: begin rd_data <= 16'h3d5b; end
				48	: begin rd_data <= 16'h3d3f; end
				49	: begin rd_data <= 16'h3d21; end
				50	: begin rd_data <= 16'h3d03; end
				51	: begin rd_data <= 16'h3ce4; end
				52	: begin rd_data <= 16'h3cc5; end
				53	: begin rd_data <= 16'h3ca5; end
				54	: begin rd_data <= 16'h3c85; end
				55	: begin rd_data <= 16'h3c64; end
				56	: begin rd_data <= 16'h3c42; end
				57	: begin rd_data <= 16'h3c20; end
				58	: begin rd_data <= 16'h3bfd; end
				59	: begin rd_data <= 16'h3bda; end
				60	: begin rd_data <= 16'h3bb6; end
				61	: begin rd_data <= 16'h3b92; end
				62	: begin rd_data <= 16'h3b6d; end
				63	: begin rd_data <= 16'h3b47; end
				64	: begin rd_data <= 16'h3b21; end
				65	: begin rd_data <= 16'h3afa; end
				66	: begin rd_data <= 16'h3ad3; end
				67	: begin rd_data <= 16'h3aab; end
				68	: begin rd_data <= 16'h3a82; end
				69	: begin rd_data <= 16'h3a59; end
				70	: begin rd_data <= 16'h3a30; end
				71	: begin rd_data <= 16'h3a06; end
				72	: begin rd_data <= 16'h39db; end
				73	: begin rd_data <= 16'h39b0; end
				74	: begin rd_data <= 16'h3984; end
				75	: begin rd_data <= 16'h3958; end
				76	: begin rd_data <= 16'h392b; end
				77	: begin rd_data <= 16'h38fd; end
				78	: begin rd_data <= 16'h38cf; end
				79	: begin rd_data <= 16'h38a1; end
				80	: begin rd_data <= 16'h3871; end
				81	: begin rd_data <= 16'h3842; end
				82	: begin rd_data <= 16'h3812; end
				83	: begin rd_data <= 16'h37e1; end
				84	: begin rd_data <= 16'h37b0; end
				85	: begin rd_data <= 16'h377e; end
				86	: begin rd_data <= 16'h374b; end
				87	: begin rd_data <= 16'h3718; end
				88	: begin rd_data <= 16'h36e5; end
				89	: begin rd_data <= 16'h36b1; end
				90	: begin rd_data <= 16'h367d; end
				91	: begin rd_data <= 16'h3648; end
				92	: begin rd_data <= 16'h3612; end
				93	: begin rd_data <= 16'h35dc; end
				94	: begin rd_data <= 16'h35a5; end
				95	: begin rd_data <= 16'h356e; end
				96	: begin rd_data <= 16'h3537; end
				97	: begin rd_data <= 16'h34ff; end
				98	: begin rd_data <= 16'h34c6; end
				99	: begin rd_data <= 16'h348d; end
				100	: begin rd_data <= 16'h3453; end
				101	: begin rd_data <= 16'h3419; end
				102	: begin rd_data <= 16'h33df; end
				103	: begin rd_data <= 16'h33a3; end
				104	: begin rd_data <= 16'h3368; end
				105	: begin rd_data <= 16'h332c; end
				106	: begin rd_data <= 16'h32ef; end
				107	: begin rd_data <= 16'h32b2; end
				108	: begin rd_data <= 16'h3274; end
				109	: begin rd_data <= 16'h3236; end
				110	: begin rd_data <= 16'h31f8; end
				111	: begin rd_data <= 16'h31b9; end
				112	: begin rd_data <= 16'h3179; end
				113	: begin rd_data <= 16'h3139; end
				114	: begin rd_data <= 16'h30f9; end
				115	: begin rd_data <= 16'h30b8; end
				116	: begin rd_data <= 16'h3076; end
				117	: begin rd_data <= 16'h3034; end
				118	: begin rd_data <= 16'h2ff2; end
				119	: begin rd_data <= 16'h2faf; end
				120	: begin rd_data <= 16'h2f6c; end
				121	: begin rd_data <= 16'h2f28; end
				122	: begin rd_data <= 16'h2ee4; end
				123	: begin rd_data <= 16'h2e9f; end
				124	: begin rd_data <= 16'h2e5a; end
				125	: begin rd_data <= 16'h2e15; end
				126	: begin rd_data <= 16'h2dcf; end
				127	: begin rd_data <= 16'h2d88; end
				128	: begin rd_data <= 16'h2d41; end
				129	: begin rd_data <= 16'h2cfa; end
				130	: begin rd_data <= 16'h2cb2; end
				131	: begin rd_data <= 16'h2c6a; end
				132	: begin rd_data <= 16'h2c21; end
				133	: begin rd_data <= 16'h2bd8; end
				134	: begin rd_data <= 16'h2b8f; end
				135	: begin rd_data <= 16'h2b45; end
				136	: begin rd_data <= 16'h2afb; end
				137	: begin rd_data <= 16'h2ab0; end
				138	: begin rd_data <= 16'h2a65; end
				139	: begin rd_data <= 16'h2a1a; end
				140	: begin rd_data <= 16'h29ce; end
				141	: begin rd_data <= 16'h2981; end
				142	: begin rd_data <= 16'h2935; end
				143	: begin rd_data <= 16'h28e7; end
				144	: begin rd_data <= 16'h289a; end
				145	: begin rd_data <= 16'h284c; end
				146	: begin rd_data <= 16'h27fe; end
				147	: begin rd_data <= 16'h27af; end
				148	: begin rd_data <= 16'h2760; end
				149	: begin rd_data <= 16'h2711; end
				150	: begin rd_data <= 16'h26c1; end
				151	: begin rd_data <= 16'h2671; end
				152	: begin rd_data <= 16'h2620; end
				153	: begin rd_data <= 16'h25cf; end
				154	: begin rd_data <= 16'h257e; end
				155	: begin rd_data <= 16'h252c; end
				156	: begin rd_data <= 16'h24da; end
				157	: begin rd_data <= 16'h2488; end
				158	: begin rd_data <= 16'h2435; end
				159	: begin rd_data <= 16'h23e2; end
				160	: begin rd_data <= 16'h238e; end
				161	: begin rd_data <= 16'h233b; end
				162	: begin rd_data <= 16'h22e7; end
				163	: begin rd_data <= 16'h2292; end
				164	: begin rd_data <= 16'h223d; end
				165	: begin rd_data <= 16'h21e8; end
				166	: begin rd_data <= 16'h2193; end
				167	: begin rd_data <= 16'h213d; end
				168	: begin rd_data <= 16'h20e7; end
				169	: begin rd_data <= 16'h2091; end
				170	: begin rd_data <= 16'h203a; end
				171	: begin rd_data <= 16'h1fe3; end
				172	: begin rd_data <= 16'h1f8c; end
				173	: begin rd_data <= 16'h1f34; end
				174	: begin rd_data <= 16'h1edc; end
				175	: begin rd_data <= 16'h1e84; end
				176	: begin rd_data <= 16'h1e2b; end
				177	: begin rd_data <= 16'h1dd3; end
				178	: begin rd_data <= 16'h1d79; end
				179	: begin rd_data <= 16'h1d20; end
				180	: begin rd_data <= 16'h1cc6; end
				181	: begin rd_data <= 16'h1c6c; end
				182	: begin rd_data <= 16'h1c12; end
				183	: begin rd_data <= 16'h1bb8; end
				184	: begin rd_data <= 16'h1b5d; end
				185	: begin rd_data <= 16'h1b02; end
				186	: begin rd_data <= 16'h1aa7; end
				187	: begin rd_data <= 16'h1a4b; end
				188	: begin rd_data <= 16'h19ef; end
				189	: begin rd_data <= 16'h1993; end
				190	: begin rd_data <= 16'h1937; end
				191	: begin rd_data <= 16'h18db; end
				192	: begin rd_data <= 16'h187e; end
				193	: begin rd_data <= 16'h1821; end
				194	: begin rd_data <= 16'h17c4; end
				195	: begin rd_data <= 16'h1766; end
				196	: begin rd_data <= 16'h1709; end
				197	: begin rd_data <= 16'h16ab; end
				198	: begin rd_data <= 16'h164c; end
				199	: begin rd_data <= 16'h15ee; end
				200	: begin rd_data <= 16'h1590; end
				201	: begin rd_data <= 16'h1531; end
				202	: begin rd_data <= 16'h14d2; end
				203	: begin rd_data <= 16'h1473; end
				204	: begin rd_data <= 16'h1413; end
				205	: begin rd_data <= 16'h13b4; end
				206	: begin rd_data <= 16'h1354; end
				207	: begin rd_data <= 16'h12f4; end
				208	: begin rd_data <= 16'h1294; end
				209	: begin rd_data <= 16'h1234; end
				210	: begin rd_data <= 16'h11d3; end
				211	: begin rd_data <= 16'h1173; end
				212	: begin rd_data <= 16'h1112; end
				213	: begin rd_data <= 16'h10b1; end
				214	: begin rd_data <= 16'h1050; end
				215	: begin rd_data <= 16'h0fee; end
				216	: begin rd_data <= 16'h0f8d; end
				217	: begin rd_data <= 16'h0f2b; end
				218	: begin rd_data <= 16'h0eca; end
				219	: begin rd_data <= 16'h0e68; end
				220	: begin rd_data <= 16'h0e06; end
				221	: begin rd_data <= 16'h0da4; end
				222	: begin rd_data <= 16'h0d41; end
				223	: begin rd_data <= 16'h0cdf; end
				224	: begin rd_data <= 16'h0c7c; end
				225	: begin rd_data <= 16'h0c1a; end
				226	: begin rd_data <= 16'h0bb7; end
				227	: begin rd_data <= 16'h0b54; end
				228	: begin rd_data <= 16'h0af1; end
				229	: begin rd_data <= 16'h0a8e; end
				230	: begin rd_data <= 16'h0a2b; end
				231	: begin rd_data <= 16'h09c7; end
				232	: begin rd_data <= 16'h0964; end
				233	: begin rd_data <= 16'h0901; end
				234	: begin rd_data <= 16'h089d; end
				235	: begin rd_data <= 16'h0839; end
				236	: begin rd_data <= 16'h07d6; end
				237	: begin rd_data <= 16'h0772; end
				238	: begin rd_data <= 16'h070e; end
				239	: begin rd_data <= 16'h06aa; end
				240	: begin rd_data <= 16'h0646; end
				241	: begin rd_data <= 16'h05e2; end
				242	: begin rd_data <= 16'h057e; end
				243	: begin rd_data <= 16'h051a; end
				244	: begin rd_data <= 16'h04b5; end
				245	: begin rd_data <= 16'h0451; end
				246	: begin rd_data <= 16'h03ed; end
				247	: begin rd_data <= 16'h0388; end
				248	: begin rd_data <= 16'h0324; end
				249	: begin rd_data <= 16'h02c0; end
				250	: begin rd_data <= 16'h025b; end
				251	: begin rd_data <= 16'h01f7; end
				252	: begin rd_data <= 16'h0192; end
				253	: begin rd_data <= 16'h012e; end
				254	: begin rd_data <= 16'h00c9; end
				255	: begin rd_data <= 16'h0065; end
				256	: begin rd_data <= 16'h0000; end
				257	: begin rd_data <= 16'hff9b; end
				258	: begin rd_data <= 16'hff37; end
				259	: begin rd_data <= 16'hfed2; end
				260	: begin rd_data <= 16'hfe6e; end
				261	: begin rd_data <= 16'hfe09; end
				262	: begin rd_data <= 16'hfda5; end
				263	: begin rd_data <= 16'hfd40; end
				264	: begin rd_data <= 16'hfcdc; end
				265	: begin rd_data <= 16'hfc78; end
				266	: begin rd_data <= 16'hfc13; end
				267	: begin rd_data <= 16'hfbaf; end
				268	: begin rd_data <= 16'hfb4b; end
				269	: begin rd_data <= 16'hfae6; end
				270	: begin rd_data <= 16'hfa82; end
				271	: begin rd_data <= 16'hfa1e; end
				272	: begin rd_data <= 16'hf9ba; end
				273	: begin rd_data <= 16'hf956; end
				274	: begin rd_data <= 16'hf8f2; end
				275	: begin rd_data <= 16'hf88e; end
				276	: begin rd_data <= 16'hf82a; end
				277	: begin rd_data <= 16'hf7c7; end
				278	: begin rd_data <= 16'hf763; end
				279	: begin rd_data <= 16'hf6ff; end
				280	: begin rd_data <= 16'hf69c; end
				281	: begin rd_data <= 16'hf639; end
				282	: begin rd_data <= 16'hf5d5; end
				283	: begin rd_data <= 16'hf572; end
				284	: begin rd_data <= 16'hf50f; end
				285	: begin rd_data <= 16'hf4ac; end
				286	: begin rd_data <= 16'hf449; end
				287	: begin rd_data <= 16'hf3e6; end
				288	: begin rd_data <= 16'hf384; end
				289	: begin rd_data <= 16'hf321; end
				290	: begin rd_data <= 16'hf2bf; end
				291	: begin rd_data <= 16'hf25c; end
				292	: begin rd_data <= 16'hf1fa; end
				293	: begin rd_data <= 16'hf198; end
				294	: begin rd_data <= 16'hf136; end
				295	: begin rd_data <= 16'hf0d5; end
				296	: begin rd_data <= 16'hf073; end
				297	: begin rd_data <= 16'hf012; end
				298	: begin rd_data <= 16'hefb0; end
				299	: begin rd_data <= 16'hef4f; end
				300	: begin rd_data <= 16'heeee; end
				301	: begin rd_data <= 16'hee8d; end
				302	: begin rd_data <= 16'hee2d; end
				303	: begin rd_data <= 16'hedcc; end
				304	: begin rd_data <= 16'hed6c; end
				305	: begin rd_data <= 16'hed0c; end
				306	: begin rd_data <= 16'hecac; end
				307	: begin rd_data <= 16'hec4c; end
				308	: begin rd_data <= 16'hebed; end
				309	: begin rd_data <= 16'heb8d; end
				310	: begin rd_data <= 16'heb2e; end
				311	: begin rd_data <= 16'heacf; end
				312	: begin rd_data <= 16'hea70; end
				313	: begin rd_data <= 16'hea12; end
				314	: begin rd_data <= 16'he9b4; end
				315	: begin rd_data <= 16'he955; end
				316	: begin rd_data <= 16'he8f7; end
				317	: begin rd_data <= 16'he89a; end
				318	: begin rd_data <= 16'he83c; end
				319	: begin rd_data <= 16'he7df; end
				320	: begin rd_data <= 16'he782; end
				321	: begin rd_data <= 16'he725; end
				322	: begin rd_data <= 16'he6c9; end
				323	: begin rd_data <= 16'he66d; end
				324	: begin rd_data <= 16'he611; end
				325	: begin rd_data <= 16'he5b5; end
				326	: begin rd_data <= 16'he559; end
				327	: begin rd_data <= 16'he4fe; end
				328	: begin rd_data <= 16'he4a3; end
				329	: begin rd_data <= 16'he448; end
				330	: begin rd_data <= 16'he3ee; end
				331	: begin rd_data <= 16'he394; end
				332	: begin rd_data <= 16'he33a; end
				333	: begin rd_data <= 16'he2e0; end
				334	: begin rd_data <= 16'he287; end
				335	: begin rd_data <= 16'he22d; end
				336	: begin rd_data <= 16'he1d5; end
				337	: begin rd_data <= 16'he17c; end
				338	: begin rd_data <= 16'he124; end
				339	: begin rd_data <= 16'he0cc; end
				340	: begin rd_data <= 16'he074; end
				341	: begin rd_data <= 16'he01d; end
				342	: begin rd_data <= 16'hdfc6; end
				343	: begin rd_data <= 16'hdf6f; end
				344	: begin rd_data <= 16'hdf19; end
				345	: begin rd_data <= 16'hdec3; end
				346	: begin rd_data <= 16'hde6d; end
				347	: begin rd_data <= 16'hde18; end
				348	: begin rd_data <= 16'hddc3; end
				349	: begin rd_data <= 16'hdd6e; end
				350	: begin rd_data <= 16'hdd19; end
				351	: begin rd_data <= 16'hdcc5; end
				352	: begin rd_data <= 16'hdc72; end
				353	: begin rd_data <= 16'hdc1e; end
				354	: begin rd_data <= 16'hdbcb; end
				355	: begin rd_data <= 16'hdb78; end
				356	: begin rd_data <= 16'hdb26; end
				357	: begin rd_data <= 16'hdad4; end
				358	: begin rd_data <= 16'hda82; end
				359	: begin rd_data <= 16'hda31; end
				360	: begin rd_data <= 16'hd9e0; end
				361	: begin rd_data <= 16'hd98f; end
				362	: begin rd_data <= 16'hd93f; end
				363	: begin rd_data <= 16'hd8ef; end
				364	: begin rd_data <= 16'hd8a0; end
				365	: begin rd_data <= 16'hd851; end
				366	: begin rd_data <= 16'hd802; end
				367	: begin rd_data <= 16'hd7b4; end
				368	: begin rd_data <= 16'hd766; end
				369	: begin rd_data <= 16'hd719; end
				370	: begin rd_data <= 16'hd6cb; end
				371	: begin rd_data <= 16'hd67f; end
				372	: begin rd_data <= 16'hd632; end
				373	: begin rd_data <= 16'hd5e6; end
				374	: begin rd_data <= 16'hd59b; end
				375	: begin rd_data <= 16'hd550; end
				376	: begin rd_data <= 16'hd505; end
				377	: begin rd_data <= 16'hd4bb; end
				378	: begin rd_data <= 16'hd471; end
				379	: begin rd_data <= 16'hd428; end
				380	: begin rd_data <= 16'hd3df; end
				381	: begin rd_data <= 16'hd396; end
				382	: begin rd_data <= 16'hd34e; end
				383	: begin rd_data <= 16'hd306; end
				384	: begin rd_data <= 16'hd2bf; end
				385	: begin rd_data <= 16'hd278; end
				386	: begin rd_data <= 16'hd231; end
				387	: begin rd_data <= 16'hd1eb; end
				388	: begin rd_data <= 16'hd1a6; end
				389	: begin rd_data <= 16'hd161; end
				390	: begin rd_data <= 16'hd11c; end
				391	: begin rd_data <= 16'hd0d8; end
				392	: begin rd_data <= 16'hd094; end
				393	: begin rd_data <= 16'hd051; end
				394	: begin rd_data <= 16'hd00e; end
				395	: begin rd_data <= 16'hcfcc; end
				396	: begin rd_data <= 16'hcf8a; end
				397	: begin rd_data <= 16'hcf48; end
				398	: begin rd_data <= 16'hcf07; end
				399	: begin rd_data <= 16'hcec7; end
				400	: begin rd_data <= 16'hce87; end
				401	: begin rd_data <= 16'hce47; end
				402	: begin rd_data <= 16'hce08; end
				403	: begin rd_data <= 16'hcdca; end
				404	: begin rd_data <= 16'hcd8c; end
				405	: begin rd_data <= 16'hcd4e; end
				406	: begin rd_data <= 16'hcd11; end
				407	: begin rd_data <= 16'hccd4; end
				408	: begin rd_data <= 16'hcc98; end
				409	: begin rd_data <= 16'hcc5d; end
				410	: begin rd_data <= 16'hcc21; end
				411	: begin rd_data <= 16'hcbe7; end
				412	: begin rd_data <= 16'hcbad; end
				413	: begin rd_data <= 16'hcb73; end
				414	: begin rd_data <= 16'hcb3a; end
				415	: begin rd_data <= 16'hcb01; end
				416	: begin rd_data <= 16'hcac9; end
				417	: begin rd_data <= 16'hca92; end
				418	: begin rd_data <= 16'hca5b; end
				419	: begin rd_data <= 16'hca24; end
				420	: begin rd_data <= 16'hc9ee; end
				421	: begin rd_data <= 16'hc9b8; end
				422	: begin rd_data <= 16'hc983; end
				423	: begin rd_data <= 16'hc94f; end
				424	: begin rd_data <= 16'hc91b; end
				425	: begin rd_data <= 16'hc8e8; end
				426	: begin rd_data <= 16'hc8b5; end
				427	: begin rd_data <= 16'hc882; end
				428	: begin rd_data <= 16'hc850; end
				429	: begin rd_data <= 16'hc81f; end
				430	: begin rd_data <= 16'hc7ee; end
				431	: begin rd_data <= 16'hc7be; end
				432	: begin rd_data <= 16'hc78f; end
				433	: begin rd_data <= 16'hc75f; end
				434	: begin rd_data <= 16'hc731; end
				435	: begin rd_data <= 16'hc703; end
				436	: begin rd_data <= 16'hc6d5; end
				437	: begin rd_data <= 16'hc6a8; end
				438	: begin rd_data <= 16'hc67c; end
				439	: begin rd_data <= 16'hc650; end
				440	: begin rd_data <= 16'hc625; end
				441	: begin rd_data <= 16'hc5fa; end
				442	: begin rd_data <= 16'hc5d0; end
				443	: begin rd_data <= 16'hc5a7; end
				444	: begin rd_data <= 16'hc57e; end
				445	: begin rd_data <= 16'hc555; end
				446	: begin rd_data <= 16'hc52d; end
				447	: begin rd_data <= 16'hc506; end
				448	: begin rd_data <= 16'hc4df; end
				449	: begin rd_data <= 16'hc4b9; end
				450	: begin rd_data <= 16'hc493; end
				451	: begin rd_data <= 16'hc46e; end
				452	: begin rd_data <= 16'hc44a; end
				453	: begin rd_data <= 16'hc426; end
				454	: begin rd_data <= 16'hc403; end
				455	: begin rd_data <= 16'hc3e0; end
				456	: begin rd_data <= 16'hc3be; end
				457	: begin rd_data <= 16'hc39c; end
				458	: begin rd_data <= 16'hc37b; end
				459	: begin rd_data <= 16'hc35b; end
				460	: begin rd_data <= 16'hc33b; end
				461	: begin rd_data <= 16'hc31c; end
				462	: begin rd_data <= 16'hc2fd; end
				463	: begin rd_data <= 16'hc2df; end
				464	: begin rd_data <= 16'hc2c1; end
				465	: begin rd_data <= 16'hc2a5; end
				466	: begin rd_data <= 16'hc288; end
				467	: begin rd_data <= 16'hc26d; end
				468	: begin rd_data <= 16'hc251; end
				469	: begin rd_data <= 16'hc237; end
				470	: begin rd_data <= 16'hc21d; end
				471	: begin rd_data <= 16'hc204; end
				472	: begin rd_data <= 16'hc1eb; end
				473	: begin rd_data <= 16'hc1d3; end
				474	: begin rd_data <= 16'hc1bb; end
				475	: begin rd_data <= 16'hc1a4; end
				476	: begin rd_data <= 16'hc18e; end
				477	: begin rd_data <= 16'hc178; end
				478	: begin rd_data <= 16'hc163; end
				479	: begin rd_data <= 16'hc14f; end
				480	: begin rd_data <= 16'hc13b; end
				481	: begin rd_data <= 16'hc128; end
				482	: begin rd_data <= 16'hc115; end
				483	: begin rd_data <= 16'hc103; end
				484	: begin rd_data <= 16'hc0f1; end
				485	: begin rd_data <= 16'hc0e0; end
				486	: begin rd_data <= 16'hc0d0; end
				487	: begin rd_data <= 16'hc0c0; end
				488	: begin rd_data <= 16'hc0b1; end
				489	: begin rd_data <= 16'hc0a3; end
				490	: begin rd_data <= 16'hc095; end
				491	: begin rd_data <= 16'hc088; end
				492	: begin rd_data <= 16'hc07b; end
				493	: begin rd_data <= 16'hc06f; end
				494	: begin rd_data <= 16'hc064; end
				495	: begin rd_data <= 16'hc059; end
				496	: begin rd_data <= 16'hc04f; end
				497	: begin rd_data <= 16'hc045; end
				498	: begin rd_data <= 16'hc03c; end
				499	: begin rd_data <= 16'hc034; end
				500	: begin rd_data <= 16'hc02c; end
				501	: begin rd_data <= 16'hc025; end
				502	: begin rd_data <= 16'hc01f; end
				503	: begin rd_data <= 16'hc019; end
				504	: begin rd_data <= 16'hc014; end
				505	: begin rd_data <= 16'hc00f; end
				506	: begin rd_data <= 16'hc00b; end
				507	: begin rd_data <= 16'hc008; end
				508	: begin rd_data <= 16'hc005; end
				509	: begin rd_data <= 16'hc003; end
				510	: begin rd_data <= 16'hc001; end
				511	: begin rd_data <= 16'hc000; end
				default : begin rd_data <= 0; end
			endcase
		end
		else begin
			rd_data <= rd_data;
		end
	end
end

endmodule
